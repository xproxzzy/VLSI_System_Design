`include "FA.v"
module AS(Out, In_1, In_2, Sel);
input        [29:0] In_1;
input        [29:0] In_2;
input        Sel;
output       [30:0] Out;
wire         [29:0] c;
wire         [30:0] In_1_31;
wire         [30:0] In_2_31;
wire         [30:0] In_2_31_Sel;

assign In_1_31[29:0] = In_1[29:0];
assign In_1_31[30] = In_1[29];
assign In_2_31[29:0] = In_2[29:0];
assign In_2_31[30] = In_2[29];
assign In_2_31_Sel[0] = In_2_31[0] ^Sel;
assign In_2_31_Sel[1] = In_2_31[1] ^Sel;
assign In_2_31_Sel[2] = In_2_31[2] ^Sel;
assign In_2_31_Sel[3] = In_2_31[3] ^Sel;
assign In_2_31_Sel[4] = In_2_31[4] ^Sel;
assign In_2_31_Sel[5] = In_2_31[5] ^Sel;
assign In_2_31_Sel[6] = In_2_31[6] ^Sel;
assign In_2_31_Sel[7] = In_2_31[7] ^Sel;
assign In_2_31_Sel[8] = In_2_31[8] ^Sel;
assign In_2_31_Sel[9] = In_2_31[9] ^Sel;
assign In_2_31_Sel[10] = In_2_31[10] ^Sel;
assign In_2_31_Sel[11] = In_2_31[11] ^Sel;
assign In_2_31_Sel[12] = In_2_31[12] ^Sel;
assign In_2_31_Sel[13] = In_2_31[13] ^Sel;
assign In_2_31_Sel[14] = In_2_31[14] ^Sel;
assign In_2_31_Sel[15] = In_2_31[15] ^Sel;
assign In_2_31_Sel[16] = In_2_31[16] ^Sel;
assign In_2_31_Sel[17] = In_2_31[17] ^Sel;
assign In_2_31_Sel[18] = In_2_31[18] ^Sel;
assign In_2_31_Sel[19] = In_2_31[19] ^Sel;
assign In_2_31_Sel[20] = In_2_31[20] ^Sel;
assign In_2_31_Sel[21] = In_2_31[21] ^Sel;
assign In_2_31_Sel[22] = In_2_31[22] ^Sel;
assign In_2_31_Sel[23] = In_2_31[23] ^Sel;
assign In_2_31_Sel[24] = In_2_31[24] ^Sel;
assign In_2_31_Sel[25] = In_2_31[25] ^Sel;
assign In_2_31_Sel[26] = In_2_31[26] ^Sel;
assign In_2_31_Sel[27] = In_2_31[27] ^Sel;
assign In_2_31_Sel[28] = In_2_31[28] ^Sel;
assign In_2_31_Sel[29] = In_2_31[29] ^Sel;
assign In_2_31_Sel[30] = In_2_31[30] ^Sel;

FA FA_1(.s(Out[0]), .carry_out(c[0]), .x(In_1_31[0]), .y(In_2_31_Sel[0]), .carry_in(Sel));
FA FA_2(.s(Out[1]), .carry_out(c[1]), .x(In_1_31[1]), .y(In_2_31_Sel[1]), .carry_in(c[0]));
FA FA_3(.s(Out[2]), .carry_out(c[2]), .x(In_1_31[2]), .y(In_2_31_Sel[2]), .carry_in(c[1]));
FA FA_4(.s(Out[3]), .carry_out(c[3]), .x(In_1_31[3]), .y(In_2_31_Sel[3]), .carry_in(c[2]));
FA FA_5(.s(Out[4]), .carry_out(c[4]), .x(In_1_31[4]), .y(In_2_31_Sel[4]), .carry_in(c[3]));
FA FA_6(.s(Out[5]), .carry_out(c[5]), .x(In_1_31[5]), .y(In_2_31_Sel[5]), .carry_in(c[4]));
FA FA_7(.s(Out[6]), .carry_out(c[6]), .x(In_1_31[6]), .y(In_2_31_Sel[6]), .carry_in(c[5]));
FA FA_8(.s(Out[7]), .carry_out(c[7]), .x(In_1_31[7]), .y(In_2_31_Sel[7]), .carry_in(c[6]));
FA FA_9(.s(Out[8]), .carry_out(c[8]), .x(In_1_31[8]), .y(In_2_31_Sel[8]), .carry_in(c[7]));
FA FA_10(.s(Out[9]), .carry_out(c[9]), .x(In_1_31[9]), .y(In_2_31_Sel[9]), .carry_in(c[8]));
FA FA_11(.s(Out[10]), .carry_out(c[10]), .x(In_1_31[10]), .y(In_2_31_Sel[10]), .carry_in(c[9]));
FA FA_12(.s(Out[11]), .carry_out(c[11]), .x(In_1_31[11]), .y(In_2_31_Sel[11]), .carry_in(c[10]));
FA FA_13(.s(Out[12]), .carry_out(c[12]), .x(In_1_31[12]), .y(In_2_31_Sel[12]), .carry_in(c[11]));
FA FA_14(.s(Out[13]), .carry_out(c[13]), .x(In_1_31[13]), .y(In_2_31_Sel[13]), .carry_in(c[12]));
FA FA_15(.s(Out[14]), .carry_out(c[14]), .x(In_1_31[14]), .y(In_2_31_Sel[14]), .carry_in(c[13]));
FA FA_16(.s(Out[15]), .carry_out(c[15]), .x(In_1_31[15]), .y(In_2_31_Sel[15]), .carry_in(c[14]));
FA FA_17(.s(Out[16]), .carry_out(c[16]), .x(In_1_31[16]), .y(In_2_31_Sel[16]), .carry_in(c[15]));
FA FA_18(.s(Out[17]), .carry_out(c[17]), .x(In_1_31[17]), .y(In_2_31_Sel[17]), .carry_in(c[16]));
FA FA_19(.s(Out[18]), .carry_out(c[18]), .x(In_1_31[18]), .y(In_2_31_Sel[18]), .carry_in(c[17]));
FA FA_20(.s(Out[19]), .carry_out(c[19]), .x(In_1_31[19]), .y(In_2_31_Sel[19]), .carry_in(c[18]));
FA FA_21(.s(Out[20]), .carry_out(c[20]), .x(In_1_31[20]), .y(In_2_31_Sel[20]), .carry_in(c[19]));
FA FA_22(.s(Out[21]), .carry_out(c[21]), .x(In_1_31[21]), .y(In_2_31_Sel[21]), .carry_in(c[20]));
FA FA_23(.s(Out[22]), .carry_out(c[22]), .x(In_1_31[22]), .y(In_2_31_Sel[22]), .carry_in(c[21]));
FA FA_24(.s(Out[23]), .carry_out(c[23]), .x(In_1_31[23]), .y(In_2_31_Sel[23]), .carry_in(c[22]));
FA FA_25(.s(Out[24]), .carry_out(c[24]), .x(In_1_31[24]), .y(In_2_31_Sel[24]), .carry_in(c[23]));
FA FA_26(.s(Out[25]), .carry_out(c[25]), .x(In_1_31[25]), .y(In_2_31_Sel[25]), .carry_in(c[24]));
FA FA_27(.s(Out[26]), .carry_out(c[26]), .x(In_1_31[26]), .y(In_2_31_Sel[26]), .carry_in(c[25]));
FA FA_28(.s(Out[27]), .carry_out(c[27]), .x(In_1_31[27]), .y(In_2_31_Sel[27]), .carry_in(c[26]));
FA FA_29(.s(Out[28]), .carry_out(c[28]), .x(In_1_31[28]), .y(In_2_31_Sel[28]), .carry_in(c[27]));
FA FA_30(.s(Out[29]), .carry_out(c[29]), .x(In_1_31[29]), .y(In_2_31_Sel[29]), .carry_in(c[28]));
FA FA_31(.s(Out[30]), .carry_out(), .x(In_1_31[30]), .y(In_2_31_Sel[30]), .carry_in(c[29]));
  
endmodule